module lcd_controller(estado,D1,D2,D3,D4,D5,D6);

	input [1:0] estado;
	output reg[7:0] D1,D2,D3,D4,D5,D6;

	always @(estado)
	begin
		case(estado)
			0: begin D1 = 70; D2 = 82; D3 = 73; D4 = 79; D5 = 32; D6 = 32; end
			1: begin D1 = 78; D2 = 79; D3 = 82; D4 = 77; D5 = 65; D6 = 76; end
			2: begin D1 = 81; D2 = 85; D3 = 69; D4 = 78; D5 = 84; D6 = 69; end
		endcase
	end

endmodule
